`timescale 1ns / 1ps

module tb_mux2(

    );
    
    reg i0,i1,i2,i3,s0,s1;
    wire y;
    
    mux2 uut(i0,i1,i2,i3,s0,s1,y);
    
    initial begin
    i0=0;i1=1;i2=0;i3=1;
    s1=0;s0=0;#10
    s1=0;s0=1;#10
    s1=1;s0=0;#10
    s1=1;s0=1;#10
    $finish;
    end
endmodule
